// Author: 0716003 鄒年城  0716079	藍世堯
module Adder(
    src1_i,
    src2_i,
    sum_o
    );

//I/O ports
input  [32-1:0]  src1_i;
input  [32-1:0]	 src2_i;
output [32-1:0]	 sum_o;

//Internal Signals
reg		 [32-1:0]  sum_o;

always @(*)
	begin
		sum_o <= src1_i + src2_i;
	end

endmodule
//test
